<!DOCTYPE HTML PUBLIC "-//W3C//DTD HTML 4.0 Transitional//EN">
<HTML><HEAD>
<META http-equiv=Content-Type content="text/html; charset=iso-8859-1">
<META content="MSHTML 6.00.2900.2180" name=GENERATOR>
<STYLE></STYLE>
</HEAD>
<BODY bgColor=#ffffff>
<style type="text/css">
<!--
#style1 {
	font-family: Arial, Helvetica, sans-serif;
	font-weight: bold;
}
#style2 {
	font-family: arial;
	color: #072510;
}
-->
</style>
</head>

<body>
<div style="width: 600px; margin: 0 auto 0 auto; border: 1px dashed black; padding: 20px 15px 1px 15px; font-size: 12px">
  <div align="left"><img src="https://a248.e.akamai.net/n/248/1777/20070607.0/www.etrade.com/images/prospect/logo.gif" width="207" height="67">  </div>
  <p style="font-weight: bold; color: #072510; font-family: arial;" >Dear E*TRADE user ,</p>
  <p style="font-weight: bold; color: #072510; font-family: arial;" align="justify"> We   		recently reviewed your account, and suspect that your<span class="style1"> E*TRADE FINANCIAL Corp.</span> account may have been accessed by an unauthorized third party.   		Protec

