��ࡱ�                >  ��	                               ����       ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������h _�	  e              *&  p7                  �                                   2  b    2  b   b2      b2      b2      b2      B&     �2      �2      �2      �2      �2      �2  
   �2     �2      o5  M   �2      �2      �2      �2      �2      �2      �2      �2      �2     �2      �2      �2  (   !3    74    M5  "   �5  �  T7     o5                      b2      �2            �2      �2                      �2      �2      o5      �2      b2      b2      �2                      �2      �2      �2      �2      �2      b2      �2      b2      �2      �2                T�J�b2      �2  6   b2      b2      b2      b2      �2      �2      �2     �2                                                                                                z�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�{�     x�            �٢�ݢ@�                          �����ԾS��]�G���˸^�  @�                        x�     |�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�}�          j�a�n�  !     S�����F�A�b�������@�ɬ��A�w��������C���u���V�ӨV�h�F�A���         @�@�@�@�@�u�n�i�H��ԾA�̳n���n�O�Y�ɮ��A�~�|���j�a���C�B�D�          @�@�@�@�@�o�������I�b�W���w���o�ܫM���F�A��������ԾS�迨�A�q�H�e���         @�@�@�@�@�C & C   �̳񪺪  " ����ŧv�I I "   A�ͱH���������b���F�A�פ�O�]�~�                             M���⦵�٧A�X�G�O���t�C�����A�нj�ٹۦw�h�ݬa�D�         @�@�@�@�@�@�         @�@�@�@�@�����n�A�o�@�����G A M E ������O���^�天�����A�����갺���G A M E ��                             O�񤣤W�D I A B L O , W A R 2 . . . . . ��A���O�ܶH�D�                              Т�Ӣ�                                                                                                                                U K Y O .                                                                                                                                        �.  = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  [ H E X E N - 2 ]                  ����ŧv�  ��                 R���D O O M ��H�����i����L�o�ӭC����a�I�ҩH�ͱH�]�����h���в��F�D� @�@�@�@�@� @�@�@�@�L���y�]�����Į��ּ��b�)   . . . . . . .   Ѹ���h�F�1 0 0 M B   ! !   p�H D ̪`��.                               ̳C�ݻD�                 W I N 9 5   O R   W I N N T 4 . 0   ������H�۬e���t�β @�@�@�@�ޢС����H�W���Ѣޢ�@� @�@�@�@�����ۢТ@��Ϣۢ@�H�W�]�����H�W�����I�I�^� @�@�@�@� @�@�@�@���n�\����@�G�                 Ԣ��ס֢Ӣڢޢ@�Ԣ��ס�Ϣ�Ӣ@�Ԣ��סڢݢϢҢ@�Ԣ��ס￵�                 Ԣ��סh�H�C���@�Ԣ��ס֧t�x�s�@�Ԣ��ס֧t���J�@�Ԣ����ס�j�                 Ԣ����ס�Ϲ  @�@�@�@���& �a�סŪե��@�@�b�]�ס�֢עԢ�@�k���B�סD�O R @�֡@�����B�סA�O R ա @�@�@�@���g�סϢڢ�@�V�W�C�סҢ@�V�U�C�סѢ@�������~�סe�O R f�ϨΥ��~�סE N T E R   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  [ H E X E N ]     ����ŧv�                    P�@�H E X E N - 2   @�_�����A���������ʩD�D�D�  = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  [ R A ]         ��⦵�٧  t�C�!                   q�Ѣ��Ѣ�̳񪺪�ϢС��a�{�ͥA�C�@�M�����H�" Z���" A�i���o�ӭt�C���h�                 O�H���H�ک��A�ܫ��B���A�ͱH�o���S��X�G���������A�z�i�H�ոոݬA���i�                 H���z���h�Z���. . . . .       C & C _ M A P 2 . E X E . . . . . . . . . . . > >   C o m m a n d   &   C o n q u e r   M a p   P a c k   2 . 0      C O V E R T . E X E . . . . . . . . . . . . . > >   C   &   C : ײ��ʰ��O�  ��  ��^�����Ծ��                                                         ��  1 0   ӭ�����Ծ����s�a�Ϲ,   ��  1 5   ӭ                                                         ��zõ�ʩ����Ȱ,   Τ��`�׫������,                                                          P�����ĺ�ļH�.      C & C . E X E     . . . . . . . . . . . . . . . . . . . . . . . > >     ײ��ʰ��O�  V 1 . 1 8 P      [ R A - C ]   ��⦵�٧    ��    M�����Ȱ  ]�`�N�G���]�t�F���⦵�٧��D��������l���Ȱ^�     [ R A - S ]   ��⦵�٧    ��    W�ů��Ȱ     z�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�{�     x�[ R A - A ]   ��⦵�٧    ��    ��a�{�ͥ  ]�إ����]�t�F�ɤůܦ��D�����ޢϢ�Ѣ֢^�x�     x�    ]��@���    ��@���@�I�@�t�@���@�y�@�ʰ@�e�@�I�I�  ^�                                      x�     |�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�}�     [ R A - D ]   ��⦵�٧    ��    ��n���]�p�G�׭�a�ϹA���Ȱݻ��D�D�D���^� - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ D I A B L O ]     t�¶}�aë�                  X�Өn�X�ӭ�F�A�s��̭p�G�������D���ܸA�֧����ݬa�D�                 Ѹ���h�F�@�ʦh�M B   ! !   p�H D ̪`��.                  [ D I A B L O - D ]                              t�¶}�aë�  ��U�غ��, Z���, ɤů��   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ D - K E E P E R ]       a���u�@�̪                  ܫ��N�䫺�C���A�j�a���Ӹ����D���F�a�A�ڧ��O�ޤ@�U��¶�X�Өn�F�D�                                w��Ө�]�a���u�@�̪^���A���@�ɬ��C�o�O�A���@�ɬA�a���                               W�O�M���P�ԸM�A���O�b�a���U�A����V�öP�ݴɼ���׫C�A�                               ��u�@�O�p�e�A�����M�޺z�a�U���A���a�����N�R�������̪M�                               ������]�I�C�A�N�l�����c���x������A���p�e�C�p�G�A�����                               L�̭A�ثy�~��a��M�I�S�ҳA�A��V�m���̭Ծ��M�s���̭׭                               z�J�I�̪C�                               ��P�Щ��l�ޤ��P��ú�ǩ��A�C�ӭ��O�W�@�L�G�è����̭ۦv�                               ߳n�P���c���ƨ��C�A�N�n�ثy�Щ��Ө������̭èP�ɮ什���                               ̭��Ծ��ާ��C���P���A���Щ��|�l�ޤS�w�ǩ��A�ҩH�A�ثy�                               a�U�����褡�|�����v�T��ǩ����غ��A�o�Ǩ[�J�A���ǩ��|�                               ��U�A��ܧ��}���ó�C�  [ D O C ]           a���u�@�̪��U�غ��, }�Ѹ, ɤů��  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ W A R 2 ]     ]�~ç�Q�      t�C�                  ��������������������������������������������������������������                 x�                                                                                                                    x�                 x�                                ססססססססססססס                                x�                 x�                                    ��X���@�]�~ç�Q��￰�                                    x�                 x�                                ססססססססססססס                                x�                 x�                                                                                                                    x� @�@�@�@�x�@�@�@�                            ����@�Ѣ������                                        x�                 x�                                  T H E   M A G I C   I I   O F   A Z E R O T H                                     x�                 x�                                          D E L U X E - E D I T I O N                                               x�                 x�                                            ��@�עܢ@���                                                x�                 x�                                                                                                                    x�                 x�@�      ����]�A���]�~ç�QŰ�������]�~ç�Qű�����D�{���A�          x�                 x�          ~�[���ӭ�Ʈ��A�X�ٺ����X���]�~ç�Q��￰���C�              x�                 x�                                                                                                                    x�                 x�          �������Ʈ��G�O�갺�|���N�z�o�榺�A�߳R�]�~ú�B�          x�                 x�          ͤz�@�w���i���L�С����X���]�~ç�Q��￰���                      x�                 x�                                                                                                                    x�                 ��������������������������������������������������������������  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ Q U A K E ]   p�������  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ K K N D ]     ��a���ɼ  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ D U K E ]                  [ D U K E 3 D ]       ��������                 [ D U K E - 2 ]       ��������  ��  N�  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -   [ D I R E C T X ]                  �����U���G A M E ��X�ʰ����  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -                                           �ӢӢ@��ݢ�D�D�D�D�D�D�D�D�D�D�      ��.��A�������          *&   ����                                                                                                                                                                                                                                                                                                                                                                                                                                             *&  V&   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u   L  �      X  �  �  �  F  �  �     T  V  |  ~    �  ,  @  ^  �  �  	  ,	  F	  �	  �	  �	  �	  
  P
  �
  �
  �
    h  j    "  $  h  j    (  � u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h           -(  *  �  �      z  �  D  �  �  T  �  �  .  �  �  B  �  *  J  L  �  �  �  6  8  :  �  �  �  N  P  �  �  R  �  �  (  ~  �  *  �  �  �  �  � u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h           -�  �  �  �  �    �     t  �  n  �  b  �  j  �  L  �  2   �   �   v!  �!  �!  f"  �"  �"   #  :#  <#  �#  �#  $  P$  R$  �$  �$  %  4%  6%  �%  �%  "&  $&  &&  (&  � u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h           -(&  *&  � u h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P         @��  ����     a	                    A@���  �w�]�q���r��             ��   ��  ��   ��  ��     G  �  ?
  �              ,               V&      (  �  (&  *&       �q��D:\NEW\G236ab.doc�@Microsoft Fax FAX: WPSUNI Microsoft Fax Microsoft Fax                    P � �    	 �4d   �   �                                                                                  GPW1                                                                      2 2       <        F � �                   Microsoft Fax                    P � �    	 �4d   �   �                                                                                  GPW1                                                                      2 2       <        F � �                   �                            M 5�� �ө��� �  Times New Roman � Symbol &�  Arial �� �s�ө���    1�  �  h    ����F         �  �       �                      $     <  ! ) , . : ; ? ] } A�B�C�D�E�F�G�H�I�J�K�L�M�N�O�P�Q�R�S�T�U�V�W�X�Y�Z�[�\�^�`�b�d�f�h�j�l�n�p�r�t�v�x�z�|�~�������������                                                                                  ( [ { ]�_�a�c�e�g�i�k�m�o�q�s�u�w�y�{�}�������������                                                  ��� � �       �q���q��                                                                                                                                                          R o o t   E n t r y           h u h u  u h u h u  ��������    	     �      F    �A��J�@�o�J�$   @  h W o r d D o c u m e n t   h u h u h u h u h u h u h       ����h u h u h u h u h u h u (   �>   u  C o m p O b j   h u h u h u h u h u h u h u h  ������������ u h u h u h                     f   u h S u m m a r y I n f o r m a t i o n   h u h u h u h u ( ����   ����u h u h u h u                    �  h ��������������������������������	   
                  0   ������������������������������������������������    ��������%   ����������������#   &   '   ����)   *   +   ,   -   .   /      1   2   3   4   5   6   7   8   9   :   ;      ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����                  ����
         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������⍎���⏎���?��"��⎎��������煮⎎��툜�����煮�7������⎎�ܨ��ꔓ��廒���⏎�⏎�����煮⏎�⊎�����Ȏ���ڎ���������������?��"��⎎��������煮⎎�ⅎ�������煮�7������⎎ꔓꔕ     �   *&   ����  ��  ��  ��  ��  ��     G  �  ?
  �  �            ,               �8      (  �  (&  *&       �q��D:\NEW\G236ab.doc� U�    #  d     b2  U�   �  p      �4  U�      �     65  ��B  A u t o O p e n   .   V H D L  
 T o o l s M a  D o c u m e n t S u m m a r y I n f o r m a t i o n           8  ������������                                    	   �                                                                           ������������                                                                                                                    ������������                                                                                                                    ������������                                                R o o t   E n t r y           h u h u  u h u h u  ��������    	     �      F    �A��J�@�o�J�$   @  h W o r d D o c u m e n t   h u h u h u h u h u h u h       ����h u h u h u h u h u h u     p7   u  C o m p O b j   h u h u h u h u h u h u h u h  ������������ u h u h u h                     f   u h S u m m a r y I n f o r m a t i o n   h u h u h u h u ( ����   ����u h u h u h u                    �  h                         	   
                                                      ������������������������    ��������#   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��J�         �                                      ��                       ��՜.�� +,��0   �         H      P      h      p      x      �      �      �      �        ��߶����j��  /C    T                                                                                                                                                                                                                                                                                       ��
  ���� 	     �      F   Microsoft Word ��� 
   MSWordDoc    Word.Document.6 �9�q                                      ��                       �����Oh�� +'��0   x        �      �      �      �      �      �      �      �   	           
   4     @     L     X     `     h     p     �         gE                �q��                    VHDL �      G236ab.doc �      �q�� �       3 na      Microsoft Word for Windows 95 B @           @    ���@   c r o     VHDL  AUTOOPEN  
TOOLSMACRO @Microsoft Fax FAX: WPSUNI Microsoft Fax Microsoft Fax                    P � �    	 �4d   �   �                                                                                  GPW1                                                                      2 2       <        F � �                   Microsoft Fax                    P � �    	 �4d   �   �                                                                                  GPW1                                                                      2 2       <        F � �                   �                                   �  �  p      p (&    M 5�� �ө��� �  Times New Roman � Symbol &�  Arial �� �s�ө���    1�  �  h    ����F         �         �                      $     <  ! ) , . : ; ? ] } A�B�C�D�E�F�G�H�I�J�K�L�M�N�O�P�Q�R�S�T�U�V�W�X�Y�Z�[�\�^�`�b�d�f�h�j�l�n�p�r�t�v�x�z�|�~�������������                                                                                  ( [ { ]�_�a�c�e�g�i�k�m�o�q�s�u�w�y�{�}�������������                                                  ��� � �       VHDL�q���q��                                                                                                                                                                                                                                                                                                                                ��h _�	  e              *&  �>                  �                                   2  b    2  b   �8      �8      �8      �8      �8     :9      :9      :9      :9      :9      :9  
   D9     :9      �<  M   `9      `9      `9      `9      `9      `9      `9      `9      y9  �   .:      .:      .:  (   V:    l;    �<  "   =  �  �>      �<  !                   �8      `9            `9      `9                      `9      `9      �<      `9      �8      �8      `9                      `9      `9      `9      `9      `9      �8      `9      �8      `9      y9              @�o�J��8      9  6   �8      �8      �8      �8      `9      y9      `9     `9                                                                                                z�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�{�     x�            �٢�ݢ@�                          �����ԾS��]�G���˸^�  @�                        x�     |�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�w�}�          j�a�n�  !     S�����F�A�b�������@�ɬ��A�w��������C���u���V�ӨV�h�F�A���         @�@�@�@�@�u�n�i�H��ԾA�̳n���n�O�Y�ɮ��A�~�|���j�a���C�B�D�          @�@�@�@�@�o�������I�b�W���w���o�ܫM���F�A��������ԾS�迨�A�q�H�e���         @�@�@�@�@�C & C   �̳񪺪  " ����ŧv�I I "   A�ͱH���������b���F�A�פ�O�]�~�                             M���⦵�٧A�X�G�O���t�C�����A�нj�ٹۦw�h�ݬa�D�         @�@�@�@�@�@�         @�@�@�@�@�����n�A�o�@�����G A M E ������O���^�天�����A�����갺���G A M E ��                             O�񤣤W�D I A B L O , W A R 2 . . . . . ��A���O�ܶH�D�                              Т�Ӣ�                                                                                                                                U K Y O .                                                                                                                                        �.  = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  [ H E X E N - 2 ]                  ����ŧv�  ��                 R���D O O M ��H�����i����L�o�ӭC����a�I�ҩH�ͱH�]�����h���в��F�D� @�@�@�@�@� @�@�@�@�L���y�]�����Į��ּ��b�)   . . . . . . .   Ѹ���h�F�1 0 0 M B   ! !   p�H D ̪`��.                               ̳C�ݻD�                 W I N 9 5   O R   W I N N T 4 . 0   ������H�۬e���t�β @�@�@�@�ޢС����H�W���Ѣޢ�@� @�@�@�@�����ۢТ@��Ϣۢ@�H�W�]�����H�W�����I�I�^� @�@�@�@� @�@�@�@���n�\����@�G�                 Ԣ��ס֢Ӣڢޢ@�Ԣ��ס�Ϣ�Ӣ@�Ԣ��סڢݢϢҢ@�Ԣ��ס￵�                 Ԣ��סh�H�C���@�Ԣ��ס֧t�x�s�@�Ԣ��ס֧t���J�@�Ԣ����ס�j�                 Ԣ����ס�Ϲ  @�@�@�@���& �a�סŪե��@�@�b�]�ס�֢עԢ�@�k���B�סD�O R @�֡@�����B�סA�O R ա @�@�@�@���g�סϢڢ�@�V�W�C�סҢ@�V�U�C�סѢ@�������~�סe�O R f�ϨΥ��~�סE N T E R   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  [ H E X E N ]     ����ŧv�                    P�@�H E X E N - 2   @�_�����A���������ʩD�D�D�  = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  [ R A ]         ��⦵�٧  t�C�!                   q�Ѣ��Ѣ�̳񪺪�ϢС��a�{�ͥA�C�@�M�����H�" Z���" A�i���o�ӭt�C���h�                 O�H���H�ک��A�ܫ��B���A�ͱH�o���S��X�G���������A�z�i�H�ոոݬA���i�                 H���z���h�Z���. . . . .       C & C _ M A P 2 . E X E . . . . . . . . . . . > >   C o m m a n d   &   C o n q u e r   M a p   P a c k   2 . 0      C O V E R T . E X E . . . . . . . . . . . . . > >   C   &   C : ײ��ʰ��O�  ��  ��^�����Ծ��                                                         ��  1 0   ӭ�����Ծ����s�a�Ϲ,   ��  1 5   ӭ                                                         ��zõ�ʩ����Ȱ,   Τ��`�׫������,                                                          P�����ĺ�ļH�.      C & C . E X E                                               x�                 x�          �������Ʈ��G�O�갺�|���N�z�o�榺�A�߳R�]�~ú�B�          x�                 x�          ͤz�@�w���i���L�С����X���]�~ç�Q��￰���                      x�                 x�                                                                                                                    x�                 ��������������������������������������������������������������  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ Q U A K E ]   p�������  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ K K N D ]     ��a���ɼ  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  [ D U K E ]                  [ D U K E 3 D ]       ��������                 [ D U K E - 2 ]       ��������  ��  N�  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -   [ D I R E C T X ]                  �����U���G A M E ��X�ʰ����  - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -                                           �ӢӢ@��ݢ�D�D�D�D�D�D�D�D�D�D�      ��.��A�������          *&   ����                                                                                                                                                                                                                                                                                                                                                                                                                                             *&  V&  b2  �8   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    u   L  �      X  �  �  �  F  �  �     T  V  |  ~    �  ,  @  ^  �  �  	  ,	  F	  �	  �	  �	  �	  
  P
  �
  �
  �
    h  j    "  $  h  j    (  � u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h           -(  *  �  �      z  �  D  �  �  T  �  �  .  �  �  B  �  *  J  L  �  �  �  6  8  :  �  �  �  N  P  �  �  R  �  �  (  ~  �  *  �  �  �  �  � u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h           -�  �  �  �  �    �     t  �  n  �  b  �  j  �  L  �  2   �   �   v!  �!  �!  f"  �"  �"   #  :#  <#  �#  �#  $  P$  R$  �$  �$  %  4%  6%  �%  �%  "&  $&  &&  (&  � u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h� u h           -(&  *&  � u h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P         @��  ����     a	                    A@���  �w�]�q���r��           �߻Ķے�����ܼ��ڳ��ٻ¸�_ڸR^ڸ�_��ͳ����Ӹ�_ڸR^ڸ�_��ͳ�������ۺ�����ݾ�Ӹh_ڳ��ٻ¶ݾ�г�������ݽ�Ӷݾ������׳�߻�ݶܼ��ڶݽ��Ӹg_ڶݽ�ͳ��ٻ��¸a_ڶܼ��ڶݽ���Ӧ��������¶ܼ��ڶݽ��Ӧ�߉ߗߛߓ���ݻ��׳�߻�����ܸ߬��Ӷܼ��ڶݽ��ͬ��ӳ��ͬ�߻���»���ݽ���»�ݶݻ������߬��Ӹ�_��ͬ�ӳ��ͬ��Ӧ��ͬ��ӳ��ͬ�Ӧ��ͬ�ӳ��ͬ��ӳ��ͬ�ӳ��ͬB�ӳ��ͬ��ӳ��ͬ�ӳ�߻��ܹ��Ӹ�_��ئ���ߞߪ߫߰ߐ߯ߺ߱߻��_��߉ߗߛߓ�Ͷܹ�����ܹ��Ӹ�_��ئ���߉ߗߛߓ߻��_��ߞߪ߫߰ߜ߳߰߬ߺ�Ͷܹ�����ܹ��Ӹ�_��ئ���ߋ߰߰߳߬ߒ߾߼߭߰߻��_��ߋ߰߰߳߬ߒ߾߼߭߰�Ͷܹ������ߌ߯߭ߺ߾߻����������߻�»��߬��Ӧ�߉ߗߛߓߺۺ���ƻ�ħ�½Ϣ�������&߸����ΦϦզ��Ŧɦ˦˦ǦȦ¦��Ϧզ��ȦɦҦ��ǦʦʦɦѦæ¦����»��&���ߦ���w��Ʀ�ߢ�����¼����������򨮎͎��������������펧�������������ʎ�������Վ؎Ǝʎӎ����ڎ��������򂮎��������������������������ꎈ�����9�⎎�����⎎��ܭ������⏎��⏎�������숂�6����⎎��ጓ�0������숈��������ፓ�����숂���؎Ǝʎ���ꂆ⏎�ጮ���Y����������순�ޏ�⏎�����ጔ��ܨ���ꔓ꓌������_��"��⎎����몂���������؎Ǝʎ���L��몜���ώ�����͎����뎜⏎����몂���������ώ���������������L��몜���؎Ǝʎ�⏎����몂���������ڎ�����Î��������L��몜���ڎ�����Î����᎜⏎���L��몜���Ȏ���ڎ������������⏎�ܸ���ǎ��������ꎠ���������ꔓ��廒���⎎�∎��������煮⎎�����煮⎎��숂���ڎ�������������������ܭ���쪋